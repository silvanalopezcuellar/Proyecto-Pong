library verilog;
use verilog.vl_types.all;
entity vga_sync_vlg_vec_tst is
end vga_sync_vlg_vec_tst;
